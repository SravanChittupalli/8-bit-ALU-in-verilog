module not_gate8
(
	input [7:0] a8,
	output [7:0] y8
);

	not_gate4 n03(a8[3:0], y8[3:0]);
	not_gate4 n47(a8[7:4], y8[7:4]);

endmodule
